** Profile: "TPS55289 Startup-Startup"  [ C:\Workspace\Bryce_Xun\Simulation\PSpice\Bryce\TPS55289\TPS55289\Release\TPS55289-PSpiceFiles\TPS55289 Startup\Startup.sim ] 

** Creating circuit file "Startup.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../generic_blocks.lib" 
.LIB "../../../tps55289.lib" 
* From [PSPICE NETLIST] section of C:\Users\a0497752\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5ms 0 20n 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\TPS55289 Startup.net" 


.END
